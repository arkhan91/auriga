module spi_slave (
    input logic spi_clk,
    input logic cs_n,
    input logic rst_n,
    input logic mosi,
    input logic miso,
    
    input logic [7:0] data_i,
    output logic [7:0] data_o
);




/// Serial to Parallel 

    
endmodule