module controller #(
    parameters
)(
    
);
    

// forwarding
endmodule : controller