//  Package: core_pkg
//
package core_pkg;
    //  Group: Typedefs
    
/////////////
// Opcodes //
/////////////

    typedef enum logic [6:0] {
        OPCODE_LOAD     = 7'b000_0000,
        OPCODE_LOAD_FP  = 7'b000_0011,
        OPCODE_MISC_MEM = 7'b000_1111,
        OPCODE_OP_IMM   = 7'b001_0011,
        OPCODE_AUIPC    = 7'b001_0111,
        OPCODE_STORE    = 7'b010_0011,
        OPCODE_OP       = 7'b011_0011,
        OPCODE_LUI      = 7'b011_0111,
        OPCODE_BRANCH   = 7'b110_0011,
        OPCODE_JALR     = 7'b110_0111,
        OPCODE_JAL      = 7'b110_1111,
        OPCODE_SYSTEM   = 7'b111_0011
      } opcode_e;
      
    //  Group: Parameters
    typedef struct packed {
        logic [4:0] rs0_addr;
        logic [4:0] rs1_addr;
        logic [4:0] rd_addr;
    } regfile_op;
    
    typedef struct packed {
        logic [11:0] imm12;
        logic [4:0]  rs1_addr;
        logic [2:0]  funct3;
        logic [4:0]  rd_addr;
        logic [6:0]  opcode;
    } Itype_inst_t;

    typedef struct packed {
        logic [6:0] imm12_5;
        logic [4:0] rs2_addr;
        logic [4:0] rs1_addr;
        logic [2:0] funct3;
        logic [6:0] imm4_0;
        logic [6:0] opcode;
    } Rtype_inst_t;

    typedef struct packed {
        logic [6:0] imm12_5;
        logic [4:0] rs2_addr;
        logic [4:0] rs1_addr;
        logic [2:0] funct3;
        logic [6:0] imm4_0;
        logic [6:0] opcode;
    } Stype_inst_t;

    typedef struct packed {
        logic [6:0] funct7;
        logic [4:0] rs2_addr;
        logic [4:0] rs1_addr;
        logic [2:0] funct3;
        logic [4:0] rd_addr;
        logic [6:0] opcode;
    } Btype_inst_t;
 
    typedef struct packed {
        logic [6:0] funct7;
        logic [4:0] rs2_addr;
        logic [4:0] rs1_addr;
        logic [2:0] funct3;
        logic [4:0] rd_addr;
        logic [6:0] opcode;
    } Jtype_inst_t;

    typedef enum logic [2:0] {
        ADD  = 3'b000,
        SLL  = 3'b001,
        SLT  = 3'b010,
        SLTU = 3'b011,
        XOR  = 3'b100,
        SRL  = 3'b101,
        OR   = 3'b110,
        AND  = 3'b111
    } alu_op_t;
    
    typedef enum logic [2:0] {
        ld_LB  = 3'b000,
        ld_LH  = 3'b001,
        ld_LW  = 3'b010,
        ld_LD  = 3'b011,
        ld_LBU = 3'b100,
        ld_LHU = 3'b101,
        ld_LWU = 3'b110
    } ld_op_t;
    
    typedef enum logic [2:0] {
        SB  = 3'b000,
        SH  = 3'b001,
        LW  = 3'b010,
        LD  = 3'b011
    } sd_op_t;
    
    typedef enum logic [2:0] {
        BEQ  = 3'b000, 
        BNE  = 3'b001, 
        BLT  = 3'b100,
        BGE  = 3'b101,
        BLTU = 3'b110,   
        BGEU = 3'b111
    } branch_op_t;

    localparam int unsigned ALU_OP_BITS = 3;
    localparam int unsigned OP_BITS = 4;


    typedef enum logic [1:0]{
        IMEM,
        REG_OPERAND,
        BYPASS
    } operand_sel_t;

    typedef struct packed {
        logic [4:0] rs1_addr;
        logic [4:0] rs2_addr;
        logic [4:0] rd_addr;
    } reg_addr_t;

    typedef struct packed {
        operand_sel_t  op_mux_sel_0;
        operand_sel_t  op_mux_sel_1;
        alu_op_t       alu_op; 
        logic          invert;
        reg_addr_t     addr;
        logic [31:0]   sign_extended;
    } core_ctrl_t;

/*
    localparam [31:0] BEQ                = 32'b?????????????????000?????1100011;
    localparam [31:0] BNE                = 32'b?????????????????001?????1100011;
    localparam [31:0] BLT                = 32'b?????????????????100?????1100011;
    localparam [31:0] BGE                = 32'b?????????????????101?????1100011;
    localparam [31:0] BLTU               = 32'b?????????????????110?????1100011;
    localparam [31:0] BGEU               = 32'b?????????????????111?????1100011;
    
    localparam [31:0] JALR               = 32'b?????????????????000?????1100111;
    localparam [31:0] JAL                = 32'b?????????????????????????1101111;
    localparam [31:0] LUI                = 32'b?????????????????????????0110111;
    localparam [31:0] AUIPC              = 32'b?????????????????????????0010111;
    
    localparam [31:0] ADDI               = 32'b?????????????????000?????0010011;
    localparam [31:0] SLLI               = 32'b000000???????????001?????0010011;
    localparam [31:0] SLTI               = 32'b?????????????????010?????0010011;
    localparam [31:0] SLTIU              = 32'b?????????????????011?????0010011;
    localparam [31:0] XORI               = 32'b?????????????????100?????0010011;
    localparam [31:0] SRLI               = 32'b000000???????????101?????0010011;
    localparam [31:0] SRAI               = 32'b010000???????????101?????0010011;
    localparam [31:0] ORI                = 32'b?????????????????110?????0010011;
    localparam [31:0] ANDI               = 32'b?????????????????111?????0010011;
    
    localparam [31:0] ADD                = 32'b0000000??????????000?????0110011;
    localparam [31:0] SUB                = 32'b0100000??????????000?????0110011;
    localparam [31:0] SLL                = 32'b0000000??????????001?????0110011;
    localparam [31:0] SLT                = 32'b0000000??????????010?????0110011;
    localparam [31:0] SLTU               = 32'b0000000??????????011?????0110011;
    localparam [31:0] XOR                = 32'b0000000??????????100?????0110011;
    localparam [31:0] SRL                = 32'b0000000??????????101?????0110011;
    localparam [31:0] SRA                = 32'b0100000??????????101?????0110011;
    localparam [31:0] OR                 = 32'b0000000??????????110?????0110011;
    localparam [31:0] AND                = 32'b0000000??????????111?????0110011;
    
    localparam [31:0] ADDIW              = 32'b?????????????????000?????0011011;
    localparam [31:0] SLLIW              = 32'b0000000??????????001?????0011011;
    localparam [31:0] SRLIW              = 32'b0000000??????????101?????0011011;
    localparam [31:0] SRAIW              = 32'b0100000??????????101?????0011011;
    
    localparam [31:0] ADDW               = 32'b0000000??????????000?????0111011;
    localparam [31:0] SUBW               = 32'b0100000??????????000?????0111011;
    localparam [31:0] SLLW               = 32'b0000000??????????001?????0111011;
    localparam [31:0] SRLW               = 32'b0000000??????????101?????0111011;
    localparam [31:0] SRAW               = 32'b0100000??????????101?????0111011;
    
    localparam [31:0] LB                 = 32'b?????????????????000?????0000011;
    localparam [31:0] LH                 = 32'b?????????????????001?????0000011;
    localparam [31:0] LW                 = 32'b?????????????????010?????0000011;
    localparam [31:0] LD                 = 32'b?????????????????011?????0000011;
    localparam [31:0] LBU                = 32'b?????????????????100?????0000011;
    localparam [31:0] LHU                = 32'b?????????????????101?????0000011;
    localparam [31:0] LWU                = 32'b?????????????????110?????0000011;
    
    localparam [31:0] SB                 = 32'b?????????????????000?????0100011;
    localparam [31:0] SH                 = 32'b?????????????????001?????0100011;
    localparam [31:0] SW                 = 32'b?????????????????010?????0100011;
    localparam [31:0] SD                 = 32'b?????????????????011?????0100011;
    
    localparam [31:0] FENCE              = 32'b?????????????????000?????0001111;
    localparam [31:0] FENCE_I            = 32'b?????????????????001?????0001111;
    localparam [31:0] MUL                = 32'b0000001??????????000?????0110011;
    localparam [31:0] MULH               = 32'b0000001??????????001?????0110011;
    localparam [31:0] MULHSU             = 32'b0000001??????????010?????0110011;
    localparam [31:0] MULHU              = 32'b0000001??????????011?????0110011;
    localparam [31:0] DIV                = 32'b0000001??????????100?????0110011;
    localparam [31:0] DIVU               = 32'b0000001??????????101?????0110011;
    localparam [31:0] REM                = 32'b0000001??????????110?????0110011;
    localparam [31:0] REMU               = 32'b0000001??????????111?????0110011;
    localparam [31:0] MULW               = 32'b0000001??????????000?????0111011;
    localparam [31:0] DIVW               = 32'b0000001??????????100?????0111011;
    localparam [31:0] DIVUW              = 32'b0000001??????????101?????0111011;
    localparam [31:0] REMW               = 32'b0000001??????????110?????0111011;
    localparam [31:0] REMUW              = 32'b0000001??????????111?????0111011;
    localparam [31:0] ANDN               = 32'b0100000??????????111?????0110011;
    localparam [31:0] ORN                = 32'b0100000??????????110?????0110011;
    localparam [31:0] XNOR               = 32'b0100000??????????100?????0110011;
    localparam [31:0] GREV               = 32'b0100000??????????001?????0110011;
    localparam [31:0] SLO                = 32'b0010000??????????001?????0110011;
    localparam [31:0] SRO                = 32'b0010000??????????101?????0110011;
    localparam [31:0] ROL                = 32'b0110000??????????001?????0110011;
    localparam [31:0] ROR                = 32'b0110000??????????101?????0110011;
    localparam [31:0] SBSET              = 32'b0010100??????????001?????0110011;
    localparam [31:0] SBCLR              = 32'b0100100??????????001?????0110011;
    localparam [31:0] SBINV              = 32'b0110100??????????001?????0110011;
    localparam [31:0] SBEXT              = 32'b0100100??????????101?????0110011;
    localparam [31:0] GREVI              = 32'b010000???????????001?????0010011;
    localparam [31:0] SLOI               = 32'b001000???????????001?????0010011;
    localparam [31:0] SROI               = 32'b001000???????????101?????0010011;
    localparam [31:0] RORI               = 32'b011000???????????101?????0010011;
    localparam [31:0] SBSETI             = 32'b001010???????????001?????0010011;
    localparam [31:0] SBCLRI             = 32'b010010???????????001?????0010011;
    localparam [31:0] SBINVI             = 32'b011010???????????001?????0010011;
    localparam [31:0] SBEXTI             = 32'b010010???????????101?????0010011;
    localparam [31:0] CMIX               = 32'b?????11??????????001?????0110011;
    localparam [31:0] CMOV               = 32'b?????11??????????101?????0110011;
    localparam [31:0] FSL                = 32'b?????10??????????001?????0110011;
    localparam [31:0] FSR                = 32'b?????10??????????101?????0110011;
    localparam [31:0] FSRI               = 32'b?????1???????????101?????0010011;
    localparam [31:0] CLZ                = 32'b011000000000?????001?????0010011;
    localparam [31:0] CTZ                = 32'b011000000001?????001?????0010011;
    localparam [31:0] PCNT               = 32'b011000000010?????001?????0010011;
    localparam [31:0] CRC32_B            = 32'b011000010000?????001?????0010011;
    localparam [31:0] CRC32_H            = 32'b011000010001?????001?????0010011;
    localparam [31:0] CRC32_W            = 32'b011000010010?????001?????0010011;
    localparam [31:0] CRC32C_B           = 32'b011000011000?????001?????0010011;
    localparam [31:0] CRC32C_H           = 32'b011000011001?????001?????0010011;
    localparam [31:0] CRC32C_W           = 32'b011000011010?????001?????0010011;
    localparam [31:0] CLMUL              = 32'b0000101??????????001?????0110011;
    localparam [31:0] CLMULR             = 32'b0000101??????????010?????0110011;
    localparam [31:0] CLMULH             = 32'b0000101??????????011?????0110011;
    localparam [31:0] MIN                = 32'b0000101??????????100?????0110011;
    localparam [31:0] MAX                = 32'b0000101??????????101?????0110011;
    localparam [31:0] MINU               = 32'b0000101??????????110?????0110011;
    localparam [31:0] MAXU               = 32'b0000101??????????111?????0110011;
    localparam [31:0] SHFL               = 32'b0000100??????????001?????0110011;
    localparam [31:0] UNSHFL             = 32'b0000100??????????101?????0110011;
    localparam [31:0] BDEP               = 32'b0000100??????????010?????0110011;
    localparam [31:0] BEXT               = 32'b0000100??????????110?????0110011;
    localparam [31:0] PACK               = 32'b0000100??????????100?????0110011;
    localparam [31:0] SHFLI              = 32'b000010???????????001?????0010011;
    localparam [31:0] UNSHFLI            = 32'b000010???????????101?????0010011;
    localparam [31:0] BMATFLIP           = 32'b011000000011?????001?????0010011;
    localparam [31:0] CRC32_D            = 32'b011000010011?????001?????0010011;
    localparam [31:0] CRC32C_D           = 32'b011000011011?????001?????0010011;
    localparam [31:0] BMATOR             = 32'b0000100??????????011?????0110011;
    localparam [31:0] BMATXOR            = 32'b0000100??????????111?????0110011;
    localparam [31:0] ADDIWU             = 32'b?????????????????100?????0011011;
    localparam [31:0] SLLIU_W            = 32'b000010???????????001?????0011011;
    localparam [31:0] ADDWU              = 32'b0000101??????????000?????0111011;
    localparam [31:0] SUBWU              = 32'b0100101??????????000?????0111011;
    localparam [31:0] ADDU_W             = 32'b0000100??????????000?????0111011;
    localparam [31:0] SUBU_W             = 32'b0100100??????????000?????0111011;
    localparam [31:0] GREVW              = 32'b0100000??????????001?????0111011;
    localparam [31:0] SLOW               = 32'b0010000??????????001?????0111011;
    localparam [31:0] SROW               = 32'b0010000??????????101?????0111011;
    localparam [31:0] ROLW               = 32'b0110000??????????001?????0111011;
    localparam [31:0] RORW               = 32'b0110000??????????101?????0111011;
    localparam [31:0] SBSETW             = 32'b0010100??????????001?????0111011;
    localparam [31:0] SBCLRW             = 32'b0100100??????????001?????0111011;
    localparam [31:0] SBINVW             = 32'b0110100??????????001?????0111011;
    localparam [31:0] SBEXTW             = 32'b0100100??????????101?????0111011;
    localparam [31:0] GREVIW             = 32'b0100000??????????001?????0011011;
    localparam [31:0] SLOIW              = 32'b0010000??????????001?????0011011;
    localparam [31:0] SROIW              = 32'b0010000??????????101?????0011011;
    localparam [31:0] RORIW              = 32'b0110000??????????101?????0011011;
    localparam [31:0] SBSETIW            = 32'b0010100??????????001?????0011011;
    localparam [31:0] SBCLRIW            = 32'b0100100??????????001?????0011011;
    localparam [31:0] SBINVIW            = 32'b0110100??????????001?????0011011;
    localparam [31:0] FSLW               = 32'b?????10??????????001?????0111011;
    localparam [31:0] FSRW               = 32'b?????10??????????101?????0111011;
    localparam [31:0] FSRIW              = 32'b?????10??????????101?????0011011;
    localparam [31:0] CLZW               = 32'b011000000000?????001?????0011011;
    localparam [31:0] CTZW               = 32'b011000000001?????001?????0011011;
    localparam [31:0] PCNTW              = 32'b011000000010?????001?????0011011;
*/
endpackage: core_pkg
