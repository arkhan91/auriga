//  Package: axi4_pkg
//
package axi4_pkg;
    //  Group: Typedefs
    typedef 
    
    //  Group: Parameters
    

    
endpackage: axi4_pkg
