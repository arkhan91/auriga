//  Package: axi4_pkg
//
package axi4_pkg;
    //  Group: Typedefs
    
    
    //  Group: Parameters
    

    
endpackage: axi4_pkg
