module mem_wb #(
    
)(
   
);
    data_memory u_data_memory();
    
endmodule : mem_wb