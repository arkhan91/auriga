module exe_mem();
    
    alu u_alu();
    mult_div u_mult_div();
endmodule : exe_mem